--------------------------------------------
-- Module Name: waveform_generation_tb
--------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

library UNISIM;
use UNISIM.VComponents.all;

Entity waveform_generation_tb Is
end waveform_generation_tb;

Architecture behavior of waveform_generation_tb Is	
	Signal a : STD_LOGIC := '0';	
	Signal g1 : STD_LOGIC := '0';	
	Signal g2 : STD_LOGIC := '1';	
		
begin
	

Insert your code here




end behavior;